interface jk_intf;
  
  logic clk;
  logic rst_n;
  logic j;
  logic k;
  logic q;
  logic q_bar;
  
endinterface