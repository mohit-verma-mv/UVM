interface or_intf;
  
  logic a;
  logic b;
  logic c;
  
endinterface